// will have checker code